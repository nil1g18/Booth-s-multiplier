//N bit multiplier, must be greater than 2
`define N_BIT 8 